
module IntOsc8Mhz (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
